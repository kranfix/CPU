library ieee;
use ieee.std_logic_1164.all;

entity flip_flops is
end entity;

architecture ff of flip_flops is
begin
end ff;
