library ieee;
use ieee.std_logic_1164.all;

entity registros_8 is
port();
end entity;

architecture registrar of registros_8 is

end registrar;
