library ieee;
use ieee.std_logic_1164.all;

entity cpu is
port(
    -- Inputs
    
    -- Outputs
);
end entity;

architecture cetral of cpu is
    signal r,p: std_logic;
    signal B: std_logic_vector(11 downto 0);
begin
end cpu;
