library ieee;
use ieee.std_logic_1164.all;

entity temp_y_cont is
end entity;

architecture temporizar of temp_y_cont is
begin
end temporizar;
