library ieee;
use ieee.std_logic_1164.all;

entity bus_comun is
end entity;

architecture comun of bus_comun is
begin
end comun;
