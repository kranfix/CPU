library ieee;
use ieee.std_logic_1164.all;

entity sumador_log is
end entity;

architecture sumar of sumador_log is
begin
end sumar;
