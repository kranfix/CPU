library ieee;
use ieee.std_logic_1164.all;

entity acumulador is
port();
end entity;

architecture acumular of acumulador is

end acumular;