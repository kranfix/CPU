library ieee;
use ieee.std_logic_1164.all;

entity cpu is
port();
end entity;

architecture cetral of cpu is

end cpu;